magic
tech sky130A
magscale 1 2
timestamp 1769110503
<< locali >>
rect 157 1968 855 2045
rect -96 -208 96 152
rect 400 -206 600 -200
rect 1056 -206 1248 152
rect 398 -208 1248 -206
rect -96 -218 1248 -208
rect -96 -395 296 -218
rect 473 -395 1248 -218
rect -96 -398 1248 -395
rect -96 -400 603 -398
<< viali >>
rect 296 -395 473 -218
<< metal1 >>
rect 154 3872 226 3960
rect 158 440 222 3872
rect 290 680 479 3887
rect 672 3768 1125 3960
rect 933 2896 1125 3768
rect 737 2704 1125 2896
rect 933 1295 1125 2704
rect 719 1103 1125 1295
rect 288 600 480 680
rect 158 360 224 440
rect 158 60 222 360
rect 290 -218 479 600
rect 933 531 1125 1103
rect 695 339 1125 531
rect 672 40 864 120
rect 290 -395 296 -218
rect 473 -395 479 -218
rect 290 -407 479 -395
use JNWATR_NCH_4C5F0  xo0<0> ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 0 0 1 0
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo0<1>
timestamp 1740610800
transform 1 0 0 0 1 800
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo1
timestamp 1740610800
transform 1 0 0 0 1 1600
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo2<0>
timestamp 1740610800
transform 1 0 0 0 1 2400
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo2<1>
timestamp 1740610800
transform 1 0 0 0 1 3200
box -184 -128 1336 928
<< labels >>
flabel metal1 s 288 600 480 680 0 FreeSans 400 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal1 s 160 360 224 440 0 FreeSans 400 0 0 0 IBPS_5U
port 2 nsew signal bidirectional
flabel metal1 s 672 40 864 120 0 FreeSans 400 0 0 0 IBNS_20U
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1152 4000
<< end >>
